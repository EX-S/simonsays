module keyboard (CLOCK_50, CLOCK2_50, KEY, FPGA_I2C_SCLK, FPGA_I2C_SDAT, AUD_XCK, 
		AUD_DACLRCK, AUD_ADCLRCK, AUD_BCLK, AUD_ADCDAT, AUD_DACDAT, PS2_DAT, PS2_CLK);
		
	input CLOCK_50, CLOCK2_50;
	input [0:0] KEY;
	// I2C Audio/Video config interface
	output FPGA_I2C_SCLK;
	inout FPGA_I2C_SDAT;
	// Audio CODEC
	output AUD_XCK;
	input AUD_DACLRCK, AUD_ADCLRCK, AUD_BCLK;
	input AUD_ADCDAT;
	output AUD_DACDAT;
	input PS2_DAT;
	input PS2_CLK;
		
		wire [7:0] out;
		
		audiotop a0 (
		.CLOCK_50(CLOCK_50), .CLOCK2_50(CLOCK2_50), .KEY(KEY), .FPGA_I2C_SCLK(FPGA_I2C_SCLK), .FPGA_I2C_SDAT(FPGA_I2C_SDAT), .AUD_XCK(AUD_XCK), 
		.AUD_DACLRCK(AUD_DACLRCK), .AUD_ADCLRCK(AUD_ADCLRCK), .AUD_BCLK(AUD_BCLK), .AUD_ADCDAT(AUD_ADCDAT), .AUD_DACDAT(AUD_DACDAT), .SW(out));
		
		keyTest k0 (.PS2_DAT(PS2_DAT), .PS2_CLK(PS2_CLK), .CLOCK_50(CLOCK_50), .KEY(KEY), .LEDR(out));
		
endmodule

